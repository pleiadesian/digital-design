library verilog;
use verilog.vl_types.all;
entity leds_flow is
end leds_flow;
