library verilog;
use verilog.vl_types.all;
entity memory_game_sim is
end memory_game_sim;
